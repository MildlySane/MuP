module sum(s, a,b);

input a;
input b;
output s;

xor(s,a,b);



endmodule
